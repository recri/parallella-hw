//
//  HPSDR - High Performance Software Defined Radio
//
//  Hermes code. 
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation; either version 2 of the License, or
//  (at your option) any later version.
//
//  This program is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this program; if not, write to the Free Software
//  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA

module xfirromI_1024(
		     clka,
		     addra,
		     douta
		     );
   input clka;
   input [9 : 0] addra;
   output reg [17 : 0] douta;
   parameter MifFile = "no_coe_file_loaded";

   (* RAM_STYLE="BLOCK_POWER2" *)

   reg [17:0] 	       ram [1023:0];
   
   initial
      $readmemh(MifFile, ram, 0, 1023);

   always @(posedge clka) begin
      douta <= ram[addra];
   end
endmodule

